* Two-Stage OTA with Miller Compensation
* GF180MCU Process

.param ibn = 6.28e-06
.param W0 = 5.02e-06
.param W1 = 3.99e-06
.param W2 = 3.14e-07
.param W5 = 2.31e-05
.param W6 = 6.28e-06
.param L0 = 5.00e-07
.param L1 = 5.00e-07
.param L2 = 5.77e-05
.param L5 = 5.00e-07
.param L6 = 5.77e-05
.param nf0 = 2
.param nf1 = 1
.param nf2 = 1
.param nf5 = 5
.param nf6 = 2
